module processor
(
    input   logic           clk, rst,
    // output  logic   [31:0]  PC,
    // input   logic   [31:0]  Instr,
    // output  logic           MemWriteD,
    // output  logic   [31:0]  ALUResult, WriteData,
    // input   logic   [31:0]  ReadData
);

// From/To Controller signals/buses
logic           RegWriteD, MemWriteD, JumpD, BranchD, ALUSrcD, 
logic   [2:0]   ALUControlD,
logic   [1:0]   ResultSrcD, ImmSrcD, 
logic   [31:0]  InstrD,
logic           PCSrcE,
logic           JumpE, BranchE, ZeroE,

// From/To Hazard Unit signals/buses
logic           StallF,
logic           StallD, FlushD,
logic   [4:0]   Rs1D, Rs2D,
logic           FlushE, 
logic   [1:0]   ForwardAE, ForwardBE,
logic   [4:0]   Rs1E, Rs2E, RdE, 
logic           RegWriteM,
logic   [4:0]   RdM,
logic           RegWriteW,
logic   [4:0]   RdW,

// From/To Instruction Memory signals/buses
logic   [31:0]  InstrF,
logic   [31:0]  PCF,

// From/To Data Memory signals/buses
logic   [31:0]  ReadDataM,
logic   [31:0]  ALUResultM, WriteDataM,
logic           MemWriteM

controller ctrl
(
    .op             (InstrD[6:0]),
    .funct3         (InstrD[14:12]),
    .funct7b5       (InstrD[30]),
    .ZeroD          (ZeroD),
    .ResultSrcD     (ResultSrcD),
    .MemWriteD      (MemWriteD),
    .PCSrcE         (PCSrcE),
    .ALUSrcD        (ALUSrcD),
    .RegWriteD      (RegWriteD),
    .JumpD          (JumpD),
    .ImmSrcD        (ImmSrcD),
    .ALUControlD    (ALUControlD)
);

data_path dp
(
    // System signals
    .clk            (clk),
    .rst            (rst),

    // From/To Controller signals/buses 
    .RegWriteD      (RegWriteD),
    .MemWriteD      (MemWriteD),
    .JumpD          (JumpD),
    .BranchD        (BranchD),
    .ALUSrcD        (ALUSrcD),
    .ALUControlD    (ALUControlD),
    .ResultSrcD     (ResultSrcD),
    .ImmSrcD        (ImmSrcD),
    .InstrD         (InstrD),

    .PCSrcE         (PCSrcE),
    .JumpE          (JumpE),
    .BranchE        (BranchE),
    .ZeroE          (ZeroE),

    // From/To Hazard Unit signals/buses
    .StallF         (StallF),

    .StallD         (StallD),
    .FlushD         (FlushD),
    .Rs1D           (Rs1D),
    .Rs2D           (Rs2D),

    .ResultSrcEb0   (ResultSrcE[0]),
    .FlushE         (FlushE),
    .ForwardAE      (ForwardAE),
    .ForwardBE      (ForwardBE),
    .Rs1E           (Rs1E),
    .Rs2E           (Rs2E),
    .RdE            (RdE),

    .RegWriteM      (RegWriteM),
    .RdM            (RdM),

    .RegWriteW      (RegWriteW),
    .RdW            (RdW),

    // From/To Instruction Memory signals/buses
    .InstrF         (InstrF),
    .PCF            (PCF),

    // From/To Data Memory signals/buses
    .ReadDataM      (ReadDataM),
    .ALUResultM     (ALUResultM),
    .WriteDataM     (WriteDataM),
    .MemWriteM      (MemWriteM)
);

hazard_unit hu
(
    .Rs1D         (Rs1D),
    .Rs2D         (Rs2D),
    .Rs1E         (Rs1E),
    .Rs2E         (Rs2E),
    .RdE          (RdE),
    .RdM          (RdM),
    .RdW          (RdW),
    .PCSrcE       (PCSrcE),
    .ResultSrcEb0 (ResultSrcE[0]),
    .RegWriteM    (RegWriteM),
    .RegWriteW    (RegWriteW),
    
    .StallF       (StallF),
    .StallD       (StallD),
    .FlushD       (FlushD),
    .FlushE       (FlushE),
    .ForwardAE    (ForwardAE),
    .ForwardBE    (ForwardBE)
);

endmodule
